module
#(
    parameter NB_OP = 6,
    parameter NB_DATA = 8,
    parameter NB_FULL_DATA = 10,
)
(

)

endmodule